package defs;
  timeunit 1ns; timeprecision 1ps;
  `include "header/cpu_profile.svh"
  `include "header/signal_types.svh"
  `include "header/decode.svh"
  `include "header/cpu_buffer_bus.svh"
  `include "header/AXI_define.svh"

endpackage
