import defs::*;

module EX #(
    parameter XLEN = 32
) ();

endmodule
