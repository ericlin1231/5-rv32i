module MEM #(
    parameter XLEN = 32,
    parameter MEM_SZIE = 4096
) ();

endmodule
