module WB #(
    parameter XLEN = 32
) ();

endmodule
