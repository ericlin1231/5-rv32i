module top #(
    parameter WIDTH = 32,
    parameter MEM_SIZE = 4096
);


endmodule
