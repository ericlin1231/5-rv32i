package defs;

`include "header/signal_types.svh"
`include "header/cpu_profile.svh"
`include "header/decode.svh"
`include "header/cpu_buffer_bus.svh"

endpackage
