module ControlUnit #(
    parameter XLEN = 32
) (
);

endmodule
