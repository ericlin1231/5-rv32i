import defs::*;
