module ID #(
    parameter XLEN = 32
) ();

endmodule
